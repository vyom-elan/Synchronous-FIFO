

`include "fifo_base_seq.sv"
