
module fifo_bind;

endmodule
