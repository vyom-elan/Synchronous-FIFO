
// base register reg class which will be used to generate the reg map
class dv_base_reg_map extends uvm_reg_map;
  `uvm_object_utils(dv_base_reg_map)
  `uvm_object_new
endclass
