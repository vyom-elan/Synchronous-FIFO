
`include "fifo_base_vseq.sv"
`include "fifo_smoke_vseq.sv"
`include "fifo_common_vseq.sv"
`include "fifo_overflow_vseq.sv"
`include "fifo_underflow_vseq.sv"
`include "fifo_almost_full_empty_vseq.sv"
`include "fifo_back_to_back_vseq.sv"
